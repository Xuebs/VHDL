work.ted_and3(ted_arch) rtlc_no_parameters
